module vapor

interface Packable {
	pack() []byte
}