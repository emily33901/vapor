module vapor

struct ConnectedCallback {
}

struct DisconnectedCallback {
}
