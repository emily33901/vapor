module vapor

import proto


