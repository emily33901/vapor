module vapor

import rand

const (
	hardcoded_cm_list = [
		'162.254.196.84:27019',
		'162.254.196.84:27018',
		'162.254.196.83:27017',
		'162.254.196.83:27018',
		'162.254.196.83:27019',
		'162.254.196.67:27017',
		'162.254.196.67:27019',
		'162.254.196.68:27018',
		'162.254.196.68:27019',
		'162.254.196.67:27018',
		'162.254.196.68:27017',
		'162.254.196.84:27017',
		'155.133.248.36:27017',
		'155.133.248.38:27019',
		'155.133.248.36:27018',
		'155.133.248.35:27018',
		'155.133.248.36:27020',
		'155.133.248.34:27017',
		'155.133.248.39:27023',
		'155.133.248.39:27022',
		'155.133.248.37:27019',
		'155.133.248.39:27024',
		'155.133.248.37:27017',
		'155.133.248.38:27026',
		'155.133.248.34:27021',
		'155.133.248.35:27021',
		'155.133.248.34:27018',
		'155.133.248.35:27019',
		'155.133.248.36:27021',
		'155.133.248.35:27020',
		'155.133.248.38:27020',
		'155.133.248.38:27024',
		'155.133.248.38:27025',
		'155.133.248.39:27025',
		'155.133.248.38:27023',
		'155.133.248.39:27020',
		'155.133.248.37:27020',
		'155.133.248.34:27019',
		'155.133.248.39:27027',
		'155.133.248.38:27021',
		'155.133.248.38:27022',
		'155.133.248.39:27018',
		'155.133.248.39:27019',
		'155.133.248.38:27017',
		'155.133.248.38:27027',
		'155.133.248.39:27026',
		'155.133.248.39:27021',
		'155.133.248.38:27018',
		'155.133.248.36:27019',
		'155.133.248.37:27018',
		'155.133.248.35:27017',
		'155.133.248.34:27020',
		'155.133.248.39:27017',
		'155.133.248.37:27021',
		'185.25.182.76:27018',
		'185.25.182.77:27019',
		'185.25.182.77:27018',
		'185.25.182.76:27020',
		'185.25.182.77:27021',
		'185.25.182.76:27021',
		'185.25.182.76:27017',
		'185.25.182.77:27020',
		'185.25.182.76:27019',
		'185.25.182.77:27017',
		'162.254.192.87:27018',
		'162.254.192.87:27023',
		'162.254.192.101:27021',
		'162.254.192.87:27019',
		'162.254.192.109:27019',
		'162.254.192.71:27017',
		'162.254.192.108:27019',
		'162.254.192.109:27017',
		'162.254.192.71:27024',
		'162.254.192.87:27026',
		'162.254.192.87:27022',
		'162.254.192.101:27018',
		'162.254.192.100:27017',
		'162.254.192.87:27020',
		'162.254.192.87:27017',
		'162.254.192.87:27025',
		'162.254.192.71:27026',
		'162.254.192.87:27021',
		'162.254.192.87:27027',
		'162.254.192.71:27025',
		'162.254.192.101:27017',
		'162.254.192.71:27022',
		'162.254.192.109:27020',
		'162.254.192.71:27021',
		'162.254.192.100:27019',
		'162.254.192.100:27021',
		'162.254.192.108:27018',
		'162.254.192.108:27021',
		'162.254.192.109:27021',
		'162.254.192.109:27018',
		'162.254.192.101:27019',
		'162.254.192.108:27020',
		'162.254.192.108:27017',
		'162.254.192.100:27020',
		'162.254.192.71:27019',
		'162.254.192.101:27020',
	]
)

fn hardcoded_cm() string {
	return hardcoded_cm_list[rand.int_in_range(0, hardcoded_cm_list.len)]
}
