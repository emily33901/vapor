module vapor

enum Msg
{
	invalid = 0
	multi = 1
	protobuf_wrapped = 2

	// base_general = 100
	generic_reply = 100
	dest_job_failed = 113
	alert = 115
	scid_request = 120
	scid_response = 121
	job_heartbeat = 123
	hub_connect = 124
	subscribe = 126
	route_message = 127
	// remote_sys_id = 128 // removed
	// am_create_account_response = 129 // obsolete
	wg_request = 130
	wg_response = 131
	keep_alive = 132
	web_api_job_request = 133
	web_api_job_response = 134
	client_session_start = 135
	client_session_end = 136
	// client_session_update_auth_ticket = 137 // removed "renamed to ClientSessionUpdate"
	client_session_update = 137
	// stats_deprecated = 138 // removed
	ping = 139
	ping_response = 140
	stats = 141
	request_full_stats_block = 142
	load_dbo_cache_item = 143
	load_dbo_cache_item_response = 144
	invalidate_dbo_cache_items = 145
	service_method = 146
	service_method_response = 147
	client_package_versions = 148
	timestamp_request = 149
	timestamp_response = 150
	service_method_call_from_client = 151
	service_method_send_to_client = 152

	// base_shell = 200
	assign_sys_id = 200
	exit = 201
	dir_request = 202
	dir_response = 203
	zip_request = 204
	zip_response = 205
	update_record_response = 215
	update_credit_card_request = 221
	update_user_ban_response = 225
	prepare_to_exit = 226
	content_description_update = 227
	test_reset_server = 228
	universe_changed = 229
	shell_config_info_update = 230
	request_windows_event_log_entries = 233
	provide_windows_event_log_entries = 234
	shell_search_logs = 235
	shell_search_logs_response = 236
	shell_check_windows_updates = 237
	shell_check_windows_updates_response = 238
	// shell_flush_user_license_cache = 239 // removed
	test_flush_delayed_sql = 240
	test_flush_delayed_sql_response = 241
	ensure_execute_scheduled_task_test = 242
	ensure_execute_scheduled_task_response_test = 243
	update_scheduled_task_enable_state_test = 244
	update_scheduled_task_enable_state_response_test = 245
	content_description_delta_update = 246

	// base_gm = 300
	heartbeat = 300
	shell_failed = 301
	exit_shells = 307
	exit_shell = 308
	graceful_exit_shell = 309
	// notify_watchdog = 314 // removed "Value changed to 10000"
	license_processing_complete = 316
	set_test_flag = 317
	queued_emails_complete = 318
	gm_report_php_error = 319
	gmdrm_sync = 320
	physical_box_inventory = 321
	update_config_file = 322
	test_init_db = 323
	gm_write_config_to_sql = 324
	gm_load_activation_codes = 325
	gm_queue_for_fbs = 326
	gm_schema_conversion_results = 327
	// gm_schema_conversion_results_response = 328 // removed
	gm_write_shell_failure_to_sql = 329
	gm_write_stats_to_sos = 330
	gm_get_service_method_routing = 331
	gm_get_service_method_routing_response = 332
	gm_convert_user_wallets = 333
	gm_test_next_build_schema_conversion = 334
	gm_test_next_build_schema_conversion_response = 335
	expect_shell_restart = 336
	hot_fix_progress = 337

	// base_ais = 400
	// ais_refresh_content_description = 401 // removed
	ais_request_content_description = 402
	ais_update_app_info = 403
	// ais_update_package_info = 404 // removed "renamed to AISUpdatePackageCosts"
	// ais_update_package_costs = 404 // obsolete
	ais_get_package_change_number = 405
	ais_get_package_change_number_response = 406
	// ais_app_info_table_changed = 407 // removed
	// ais_update_package_costs_response = 408 // obsolete
	// ais_create_marketing_message = 409 // obsolete
	// ais_create_marketing_message_response = 410 // obsolete
	// ais_get_marketing_message = 411 // obsolete
	// ais_get_marketing_message_response = 412 // obsolete
	// ais_update_marketing_message = 413 // obsolete
	// ais_update_marketing_message_response = 414 // obsolete
	// ais_request_marketing_message_update = 415 // obsolete
	// ais_delete_marketing_message = 416 // obsolete
	// ais_get_marketing_treatments = 419 // removed
	// ais_get_marketing_treatments_response = 420 // removed
	// ais_request_marketing_treatment_update = 421 // removed
	// ais_test_add_package = 422 // removed
	ai_get_app_gc_flags = 423
	ai_get_app_gc_flags_response = 424
	ai_get_app_list = 425
	ai_get_app_list_response = 426
	// ai_get_app_info = 427 // removed
	// ai_get_app_info_response = 428 // removed
	ais_get_coupon_definition = 429
	ais_get_coupon_definition_response = 430
	ais_update_slave_content_description = 431
	ais_update_slave_content_description_response = 432
	ais_test_enable_gc = 433

	// base_am = 500
	am_update_user_ban_request = 504
	am_add_license = 505
	// am_begin_processing_licenses = 507 // removed
	am_send_system_im_to_user = 508
	am_extend_license = 509
	am_add_minutes_to_license = 510
	am_cancel_license = 511
	am_init_purchase = 512
	am_purchase_response = 513
	am_get_final_price = 514
	am_get_final_price_response = 515
	am_get_legacy_game_key = 516
	am_get_legacy_game_key_response = 517
	am_find_hung_transactions = 518
	am_set_account_trusted_request = 519
	// am_complete_purchase = 521 // obsolete
	am_cancel_purchase = 522
	am_new_challenge = 523
	am_load_oem_tickets = 524
	am_fix_pending_purchase = 525
	am_fix_pending_purchase_response = 526
	am_is_user_banned = 527
	am_register_key = 528
	am_load_activation_codes = 529
	am_load_activation_codes_response = 530
	am_lookup_key_response = 531
	am_lookup_key = 532
	am_chat_cleanup = 533
	am_clan_cleanup = 534
	am_fix_pending_refund = 535
	am_reverse_chargeback = 536
	am_reverse_chargeback_response = 537
	am_clan_cleanup_list = 538
	am_get_licenses = 539
	am_get_licenses_response = 540
	am_send_cart_repurchase = 541
	am_send_cart_repurchase_response = 542
	allow_user_to_play_query = 550
	allow_user_to_play_response = 551
	am_verfiy_user = 552
	am_client_not_playing = 553
	// client_request_friendship = 554 // obsolete "Renamed to AMClientRequestFriendship"
	am_client_request_friendship = 554
	am_relay_publish_status = 555
	// am_reset_community_content = 556 // removed
	// am_prime_persona_state_cache = 557 // removed
	// am_allow_user_content_query = 558 // removed
	// am_allow_user_content_response = 559 // removed
	am_init_purchase_response = 560
	am_revoke_purchase_response = 561
	// am_lock_profile = 562 // removed
	am_refresh_guest_passes = 563
	// am_invite_user_to_clan = 564 // obsolete
	// am_acknowledge_clan_invite = 565 // obsolete
	am_grant_guest_passes = 566
	am_clan_data_updated = 567
	am_reload_account = 568
	am_client_chat_msg_relay = 569
	am_chat_multi = 570
	am_client_chat_invite_relay = 571
	am_chat_invite = 572
	am_client_join_chat_relay = 573
	am_client_chat_member_info_relay = 574
	am_publish_chat_member_info = 575
	am_client_accept_friend_invite = 576
	am_chat_enter = 577
	am_client_publish_removal_from_source = 578
	am_chat_action_result = 579
	am_find_accounts = 580
	am_find_accounts_response = 581
	am_request_account_data = 582
	am_request_account_data_response = 583
	am_set_account_flags = 584
	am_create_clan = 586
	am_create_clan_response = 587
	am_get_clan_details = 588
	am_get_clan_details_response = 589
	am_set_persona_name = 590
	am_set_avatar = 591
	am_authenticate_user = 592
	am_authenticate_user_response = 593
	// am_get_account_friends_count = 594 // removed
	// am_get_account_friends_count_response = 595 // removed
	amp2_p_introducer_message = 596
	client_chat_action = 597
	am_client_chat_action_relay = 598

	// base_vs = 600
	req_challenge = 600
	vac_response = 601
	req_challenge_test = 602
	vs_mark_cheat = 604
	vs_add_cheat = 605
	vs_purge_code_mod_db = 606
	vs_get_challenge_results = 607
	vs_challenge_result_text = 608
	vs_report_lingerer = 609
	vs_request_managed_challenge = 610
	vs_load_db_finished = 611

	// base_drms = 625
	drm_build_blob_request = 628
	drm_build_blob_response = 629
	drm_resolve_guid_request = 630
	drm_resolve_guid_response = 631
	drm_variability_report = 633
	drm_variability_report_response = 634
	drm_stability_report = 635
	drm_stability_report_response = 636
	drm_details_report_request = 637
	drm_details_report_response = 638
	drm_process_file = 639
	drm_admin_update = 640
	drm_admin_update_response = 641
	drm_sync = 642
	drm_sync_response = 643
	drm_process_file_response = 644
	drm_empty_guid_cache = 645
	drm_empty_guid_cache_response = 646

	// base_cs = 650
	// cs_user_content_request = 652 // removed

	// base_client = 700
	// client_log_on_deprecated = 701 // removed
	// client_anon_log_on_deprecated = 702 // removed
	client_heart_beat = 703
	client_vac_response = 704
	// client_games_played_obsolete = 705 // removed
	client_log_off = 706
	client_no_udp_connectivity = 707
	// client_inform_of_create_account = 708 // obsolete
	// client_ack_vac_ban = 709 // removed
	client_connection_stats = 710
	// client_init_purchase = 711 // removed
	client_ping_response = 712
	client_remove_friend = 714
	client_games_played_no_data_blob = 715
	client_change_status = 716
	client_vac_status_response = 717
	client_friend_msg = 718
	// client_game_connect_obsolete = 719 // removed
	// client_games_played2_obsolete = 720 // removed
	// client_game_ended_obsolete = 721 // removed
	// client_get_final_price = 722 // removed
	client_system_im = 726
	client_system_im_ack = 727
	client_get_licenses = 728
	// client_cancel_license = 729 // removed
	client_get_legacy_game_key = 730
	// client_content_server_log_on_deprecated = 731 // removed
	client_ack_vac_ban2 = 732
	// client_ack_message_by_gid = 735 // removed
	client_get_purchase_receipts = 736
	// client_ack_purchase_receipt = 737 // removed
	// client_games_played3_obsolete = 738 // removed
	// client_send_guest_pass = 739 // removed
	client_ack_guest_pass = 740
	client_redeem_guest_pass = 741
	client_games_played = 742
	client_register_key = 743
	client_invite_user_to_clan = 744
	client_acknowledge_clan_invite = 745
	client_purchase_with_machine_id = 746
	client_app_usage_event = 747
	// client_get_gift_target_list = 748 // removed
	// client_get_gift_target_list_response = 749 // removed
	client_log_on_response = 751
	// client_vac_challenge = 753 // removed
	client_set_heartbeat_rate = 755
	// client_not_logged_on_deprecated = 756 // removed
	client_logged_off = 757
	gs_approve = 758
	gs_deny = 759
	gs_kick = 760
	client_create_acct_response = 761
	client_purchase_response = 763
	client_ping = 764
	client_nop = 765
	client_persona_state = 766
	client_friends_list = 767
	client_account_info = 768
	// client_vac_status_query = 770 // removed
	client_news_update = 771
	client_game_connect_deny = 773
	gs_status_reply = 774
	// client_get_final_price_response = 775 // removed
	client_game_connect_tokens = 779
	client_license_list = 780
	// client_cancel_license_response = 781 // removed
	client_vac_ban_status = 782
	client_cm_list = 783
	client_encrypt_pct = 784
	client_get_legacy_game_key_response = 785
	// client_favorites_list = 786 // removed
	// cs_user_content_approve = 787 // removed
	// cs_user_content_deny = 788 // removed
	// client_init_purchase_response = 789 // removed
	client_add_friend = 791
	client_add_friend_response = 792
	// client_invite_friend = 793 // removed
	// client_invite_friend_response = 794 // removed
	// client_send_guest_pass_response = 795 // removed
	client_ack_guest_pass_response = 796
	client_redeem_guest_pass_response = 797
	client_update_guest_passes_list = 798
	client_chat_msg = 799
	client_chat_invite = 800
	client_join_chat = 801
	client_chat_member_info = 802
	// client_log_on_with_credentials_deprecated = 803 // removed
	client_password_change_response = 805
	client_chat_enter = 807
	client_friend_removed_from_source = 808
	client_create_chat = 809
	client_create_chat_response = 810
	// client_update_chat_metadata = 811 // removed
	client_p2_p_introducer_message = 813
	client_chat_action_result = 814
	client_request_friend_data = 815
	client_get_user_stats = 818
	client_get_user_stats_response = 819
	client_store_user_stats = 820
	client_store_user_stats_response = 821
	client_clan_state = 822
	client_service_module = 830
	client_service_call = 831
	client_service_call_response = 832
	// client_package_info_request = 833 // removed
	// client_package_info_response = 834 // removed
	client_nat_traversal_stat_event = 839
	// client_app_info_request = 840 // removed
	// client_app_info_response = 841 // removed
	client_steam_usage_event = 842
	client_check_password = 845
	client_reset_password = 846
	client_check_password_response = 848
	client_reset_password_response = 849
	client_session_token = 850
	client_drm_problem_report = 851
	client_set_ignore_friend = 855
	client_set_ignore_friend_response = 856
	client_get_app_ownership_ticket = 857
	client_get_app_ownership_ticket_response = 858
	client_get_lobby_list_response = 860
	// client_get_lobby_metadata = 861 // removed
	// client_get_lobby_metadata_response = 862 // removed
	// client_vtt_cert = 863 // removed
	// client_app_info_update = 866 // removed
	// client_app_info_changes = 867 // removed
	client_server_list = 880
	client_email_change_response = 891
	client_secret_qa_change_response = 892
	client_drm_blob_request = 896
	client_drm_blob_response = 897
	// client_lookup_key = 898 // removed
	// client_lookup_key_response = 899 // removed

	// base_game_server = 900
	gs_disconnect_notice = 901
	gs_status = 903
	gs_user_playing = 905
	gs_status2 = 906
	gs_status_update_unused = 907
	gs_server_type = 908
	gs_player_list = 909
	gs_get_user_achievement_status = 910
	gs_get_user_achievement_status_response = 911
	gs_get_play_stats = 918
	gs_get_play_stats_response = 919
	gs_get_user_group_status = 920
	am_get_user_group_status = 921
	am_get_user_group_status_response = 922
	gs_get_user_group_status_response = 923
	gs_get_reputation = 936
	gs_get_reputation_response = 937
	gs_associate_with_clan = 938
	gs_associate_with_clan_response = 939
	gs_compute_new_player_compatibility = 940
	gs_compute_new_player_compatibility_response = 941

	// base_admin = 1000
	admin_cmd = 1000
	admin_cmd_response = 1004
	admin_log_listen_request = 1005
	admin_log_event = 1006
	// log_search_request = 1007 // removed
	// log_search_response = 1008 // removed
	// log_search_cancel = 1009 // removed
	universe_data = 1010
	// request_stat_history = 1014 // removed
	// stat_history = 1015 // removed
	// admin_pw_logon = 1017 // removed
	// admin_pw_logon_response = 1018 // removed
	admin_spew = 1019
	admin_console_title = 1020
	admin_gc_spew = 1023
	admin_gc_command = 1024
	admin_gc_get_command_list = 1025
	admin_gc_get_command_list_response = 1026
	fbs_connection_data = 1027
	admin_msg_spew = 1028

	// base_fbs = 1100
	fbs_req_version = 1100
	fbs_version_info = 1101
	fbs_force_refresh = 1102
	fbs_force_bounce = 1103
	fbs_deploy_package = 1104
	fbs_deploy_response = 1105
	fbs_update_bootstrapper = 1106
	fbs_set_state = 1107
	fbs_apply_os_updates = 1108
	fbs_run_cmd_script = 1109
	fbs_reboot_box = 1110
	fbs_set_big_brother_mode = 1111
	fbs_minidump_server = 1112
	// fbs_set_shell_count_obsolete = 1113 // removed
	fbs_deploy_hot_fix_package = 1114
	fbs_deploy_hot_fix_response = 1115
	fbs_download_hot_fix = 1116
	fbs_download_hot_fix_response = 1117
	fbs_update_target_config_file = 1118
	fbs_apply_account_cred = 1119
	fbs_apply_account_cred_response = 1120
	fbs_set_shell_count = 1121
	fbs_terminate_shell = 1122
	fbs_query_gm_for_request = 1123
	fbs_query_gm_response = 1124
	fbs_terminate_zombies = 1125
	fbs_info_from_bootstrapper = 1126
	fbs_reboot_box_response = 1127
	fbs_bootstrapper_package_request = 1128
	fbs_bootstrapper_package_response = 1129
	fbs_bootstrapper_get_package_chunk = 1130
	fbs_bootstrapper_get_package_chunk_response = 1131
	fbs_bootstrapper_package_transfer_progress = 1132
	fbs_restart_bootstrapper = 1133
	fbs_pause_frozen_dumps = 1134

	// base_file_xfer = 1200
	file_xfer_request = 1200
	file_xfer_response = 1201
	file_xfer_data = 1202
	file_xfer_end = 1203
	file_xfer_data_ack = 1204

	// base_channel_auth = 1300
	channel_auth_challenge = 1300
	channel_auth_response = 1301
	channel_auth_result = 1302
	channel_encrypt_request = 1303
	channel_encrypt_response = 1304
	channel_encrypt_result = 1305

	// base_bs = 1400
	bs_purchase_start = 1401
	bs_purchase_response = 1402
	bs_authenticate_cc_trans = 1403
	bs_authenticate_cc_trans_response = 1404
	// bs_settle_nova = 1404 // removed
	bs_settle_complete = 1406
	// bs_banned_request = 1407 // removed
	bs_init_pay_pal_txn = 1408
	bs_init_pay_pal_txn_response = 1409
	bs_get_pay_pal_user_info = 1410
	bs_get_pay_pal_user_info_response = 1411
	// bs_refund_txn = 1413 // removed
	// bs_refund_txn_response = 1414 // removed
	// bs_get_events = 1415 // removed
	// bs_chase_rfr_request = 1416 // removed
	bs_payment_instr_ban = 1417
	bs_payment_instr_ban_response = 1418
	// bs_process_gc_reports = 1419 // removed
	// bs_process_pp_reports = 1420 // removed
	bs_init_gc_bank_xfer_txn = 1421
	bs_init_gc_bank_xfer_txn_response = 1422
	// bs_query_gc_bank_xfer_txn = 1423 // removed
	// bs_query_gc_bank_xfer_txn_response = 1424 // removed
	bs_commit_gc_txn = 1425
	bs_query_transaction_status = 1426
	bs_query_transaction_status_response = 1427
	// bs_query_cb_order_status = 1428 // removed
	// bs_query_cb_order_status_response = 1429 // removed
	// bs_run_red_flag_report = 1430 // removed
	bs_query_payment_inst_usage = 1431
	bs_query_payment_inst_response = 1432
	bs_query_txn_extended_info = 1433
	bs_query_txn_extended_info_response = 1434
	bs_update_conversion_rates = 1435
	// bs_process_us_bank_reports = 1436 // removed
	bs_purchase_run_fraud_checks = 1437
	bs_purchase_run_fraud_checks_response = 1438
	// bs_start_shipping_jobs = 1439 // removed
	bs_query_bank_information = 1440
	bs_query_bank_information_response = 1441
	bs_validate_xsolla_signature = 1445
	bs_validate_xsolla_signature_response = 1446
	bs_qiwi_wallet_invoice = 1448
	bs_qiwi_wallet_invoice_response = 1449
	bs_update_inventory_from_pro_pack = 1450
	bs_update_inventory_from_pro_pack_response = 1451
	bs_send_shipping_request = 1452
	bs_send_shipping_request_response = 1453
	bs_get_pro_pack_order_status = 1454
	bs_get_pro_pack_order_status_response = 1455
	bs_check_job_running = 1456
	bs_check_job_running_response = 1457
	bs_reset_package_purchase_rate_limit = 1458
	bs_reset_package_purchase_rate_limit_response = 1459
	bs_update_payment_data = 1460
	bs_update_payment_data_response = 1461
	bs_get_billing_address = 1462
	bs_get_billing_address_response = 1463
	bs_get_credit_card_info = 1464
	bs_get_credit_card_info_response = 1465
	bs_remove_expired_payment_data = 1468
	bs_remove_expired_payment_data_response = 1469
	bs_convert_to_current_keys = 1470
	bs_convert_to_current_keys_response = 1471
	bs_init_purchase = 1472
	bs_init_purchase_response = 1473
	bs_complete_purchase = 1474
	bs_complete_purchase_response = 1475
	bs_prune_card_usage_stats = 1476
	bs_prune_card_usage_stats_response = 1477
	bs_store_bank_information = 1478
	bs_store_bank_information_response = 1479
	bs_verify_posa_key = 1480
	bs_verify_posa_key_response = 1481
	bs_reverse_redeem_posa_key = 1482
	bs_reverse_redeem_posa_key_response = 1483
	bs_query_find_credit_card = 1484
	bs_query_find_credit_card_response = 1485
	bs_status_inquiry_posa_key = 1486
	bs_status_inquiry_posa_key_response = 1487
	// bs_validate_mo_pay_signature = 1488 // obsolete
	// bs_validate_mo_pay_signature_response = 1489 // obsolete
	// bs_mo_pay_confirm_product_delivery = 1490 // obsolete
	// bs_mo_pay_confirm_product_delivery_response = 1491 // obsolete
	// bs_generate_mo_pay_md5 = 1492 // obsolete
	// bs_generate_mo_pay_md5_response = 1493 // obsolete
	bs_boa_compra_confirm_product_delivery = 1494
	bs_boa_compra_confirm_product_delivery_response = 1495
	bs_generate_boa_compra_md5 = 1496
	bs_generate_boa_compra_md5_response = 1497
	bs_commit_wp_txn = 1498
	bs_commit_adyen_txn = 1499

	// base_ats = 1500
	ats_start_stress_test = 1501
	ats_stop_stress_test = 1502
	ats_run_fail_server_test = 1503
	atsufs_perf_test_task = 1504
	atsufs_perf_test_response = 1505
	ats_cycle_tcm = 1506
	ats_init_drms_stress_test = 1507
	ats_call_test = 1508
	ats_call_test_reply = 1509
	ats_start_external_stress = 1510
	ats_external_stress_job_start = 1511
	ats_external_stress_job_queued = 1512
	ats_external_stress_job_running = 1513
	ats_external_stress_job_stopped = 1514
	ats_external_stress_job_stop_all = 1515
	ats_external_stress_action_result = 1516
	ats_started = 1517
	atscs_perf_test_task = 1518
	atscs_perf_test_response = 1519

	// base_dp = 1600
	dp_set_publishing_state = 1601
	// dp_game_played_stats = 1602 // removed
	dp_unique_players_stat = 1603
	dp_streaming_unique_players_stat = 1604
	// dp_vac_infraction_stats = 1605 // obsolete
	// dp_vac_ban_stats = 1606 // obsolete
	dp_blocking_stats = 1607
	dp_nat_traversal_stats = 1608
	// dp_steam_usage_event = 1609 // removed
	// dp_vac_cert_ban_stats = 1610 // obsolete
	// dp_vac_cafe_ban_stats = 1611 // obsolete
	dp_cloud_stats = 1612
	dp_achievement_stats = 1613
	// dp_account_creation_stats = 1614 // obsolete
	dp_get_player_count = 1615
	dp_get_player_count_response = 1616
	dp_game_servers_players_stats = 1617
	// dp_download_rate_statistics = 1618 // removed
	// dp_facebook_statistics = 1619 // obsolete
	client_dp_check_special_survey = 1620
	client_dp_check_special_survey_response = 1621
	client_dp_send_special_survey_response = 1622
	client_dp_send_special_survey_response_reply = 1623
	dp_store_sale_statistics = 1624
	client_dp_update_app_job_report = 1625
	// client_dp_steam2_app_started = 1627 // removed
	dp_update_content_event = 1626
	client_dp_unsigned_install_script = 1627
	dp_partner_micro_txns = 1628
	dp_partner_micro_txns_response = 1629
	client_dp_content_stats_report = 1630
	dpvr_unique_players_stat = 1631

	// base_cm = 1700
	cm_set_allow_state = 1701
	cm_spew_allow_state = 1702
	cm_session_rejected = 1703
	cm_set_secrets = 1704
	cm_get_secrets = 1705
	// cm_app_info_response_deprecated = 1703 // removed

	// // base_dss = 1800 // removed
	// dss_new_file = 1801 // removed
	// dss_current_file_list = 1802 // removed
	// dss_synch_list = 1803 // removed
	// dss_synch_list_response = 1804 // removed
	// dss_synch_subscribe = 1805 // removed
	// dss_synch_unsubscribe = 1806 // removed

	// // base_epm = 1900 // removed
	// epm_start_process = 1901 // removed
	// epm_stop_process = 1902 // removed
	// epm_restart_process = 1903 // removed

	// base_gc = 2200
	// gc_send_client = 2200 // removed
	// am_relay_to_gc = 2201 // removed
	// gc_update_played_state = 2202 // removed
	gc_cmd_revive = 2203
	// gc_cmd_bounce = 2204 // removed
	// gc_cmd_force_bounce = 2205 // removed
	gc_cmd_down = 2206
	gc_cmd_deploy = 2207
	gc_cmd_deploy_response = 2208
	gc_cmd_switch = 2209
	am_refresh_sessions = 2210
	// gc_update_gs_state = 2211 // removed
	gc_achievement_awarded = 2212
	gc_system_message = 2213
	// gc_validate_session = 2214 // removed
	// gc_validate_session_response = 2215 // removed
	gc_cmd_status = 2216
	// gc_register_web_interfaces = 2217 // removed
	// gc_register_web_interfaces_deprecated = 2217 // removed
	// gc_get_account_details = 2218 // removed
	// gc_get_account_details_deprecated = 2218 // removed
	gc_inter_app_message = 2219
	gc_get_email_template = 2220
	gc_get_email_template_response = 2221
	// is_relay_to_gch = 2222 // removed "renamed to GCHRelay"
	gch_relay = 2222
	// gch_relay_client_to_is = 2223 // removed "renamed to GCHRelayToClient"
	gch_relay_to_client = 2223
	gch_update_session = 2224
	gch_request_update_session = 2225
	gch_request_status = 2226
	gch_request_status_response = 2227
	gch_account_vac_status_change = 2228
	gch_spawn_gc = 2229
	gch_spawn_gc_response = 2230
	gch_kill_gc = 2231
	gch_kill_gc_response = 2232
	gch_account_trade_ban_status_change = 2233
	gch_account_lock_status_change = 2234
	gch_vac_verification_change = 2235
	gch_account_phone_number_change = 2236
	gch_account_two_factor_change = 2237
	gch_invite_user_to_lobby = 2238

	// base_p2_p = 2500
	p2_p_introducer_message = 2502

	// base_sm = 2900
	sm_expensive_report = 2902
	sm_hourly_report = 2903
	// sm_fishing_report = 2904 // obsolete
	sm_partition_renames = 2905
	sm_monitor_space = 2906
	sm_test_next_build_schema_conversion = 2907
	sm_test_next_build_schema_conversion_response = 2908
	// sm_get_schema_conversion_results = 2907 // removed
	// sm_get_schema_conversion_results_response = 2908 // removed

	// base_test = 3000
	fail_server = 3000
	job_heartbeat_test = 3001
	job_heartbeat_test_response = 3002

	// base_fts_range = 3100
	// fts_get_browse_counts = 3101 // removed
	// fts_get_browse_counts_response = 3102 // removed
	// fts_browse_clans = 3103 // removed
	// fts_browse_clans_response = 3104 // removed
	// fts_search_clans_by_location = 3105 // removed
	// fts_search_clans_by_location_response = 3106 // removed
	// fts_search_players_by_location = 3107 // removed
	// fts_search_players_by_location_response = 3108 // removed
	// fts_clan_deleted = 3109 // removed
	// fts_search = 3110 // removed
	// fts_search_response = 3111 // removed
	// fts_search_status = 3112 // removed
	// fts_search_status_response = 3113 // removed
	// fts_get_gs_play_stats = 3114 // removed
	// fts_get_gs_play_stats_response = 3115 // removed
	// fts_get_gs_play_stats_for_server = 3116 // removed
	// fts_get_gs_play_stats_for_server_response = 3117 // removed
	// fts_report_ip_updates = 3118 // removed

	// base_ccs_range = 3150
	// ccs_get_comments = 3151 // removed
	// ccs_get_comments_response = 3152 // removed
	// ccs_add_comment = 3153 // removed
	// ccs_add_comment_response = 3154 // removed
	// ccs_delete_comment = 3155 // removed
	// ccs_delete_comment_response = 3156 // removed
	// ccs_preload_comments = 3157 // removed
	// ccs_notify_comment_count = 3158 // removed
	// ccs_get_comments_for_news = 3159 // removed
	// ccs_get_comments_for_news_response = 3160 // removed
	ccs_delete_all_comments_by_author = 3161
	ccs_delete_all_comments_by_author_response = 3162


	// base_lbs_range = 3200
	lbs_set_score = 3201
	lbs_set_score_response = 3202
	lbs_find_or_create_lb = 3203
	lbs_find_or_create_lb_response = 3204
	lbs_get_lb_entries = 3205
	lbs_get_lb_entries_response = 3206
	lbs_get_lb_list = 3207
	lbs_get_lb_list_response = 3208
	lbs_set_lb_details = 3209
	lbs_delete_lb = 3210
	lbs_delete_lb_entry = 3211
	lbs_reset_lb = 3212
	lbs_reset_lb_response = 3213
	lbs_delete_lb_response = 3214

	// base_ogs = 3400
	ogs_begin_session = 3401
	ogs_begin_session_response = 3402
	ogs_end_session = 3403
	ogs_end_session_response = 3404
	ogs_write_app_session_row = 3406

	// base_brp = 3600
	// brp_start_shipping_jobs = 3601 // obsolete
	// brp_process_us_bank_reports = 3602 // obsolete
	// brp_process_gc_reports = 3603 // obsolete
	// brp_process_pp_reports = 3604 // obsolete
	// brp_settle_nova = 3605 // removed
	// brp_settle_cb = 3606 // removed
	// brp_commit_gc = 3607 // obsolete
	// brp_commit_gc_response = 3608 // obsolete
	// brp_find_hung_transactions = 3609 // obsolete
	// brp_check_finance_close_out_date = 3610 // obsolete
	// brp_process_licenses = 3611 // obsolete
	// brp_process_licenses_response = 3612 // obsolete
	// brp_remove_expired_payment_data = 3613 // obsolete
	// brp_remove_expired_payment_data_response = 3614 // obsolete
	// brp_convert_to_current_keys = 3615 // obsolete
	// brp_convert_to_current_keys_response = 3616 // obsolete
	// brp_prune_card_usage_stats = 3617 // obsolete
	// brp_prune_card_usage_stats_response = 3618 // obsolete
	// brp_check_activation_codes = 3619 // obsolete
	// brp_check_activation_codes_response = 3620 // obsolete
	// brp_commit_wp = 3621 // obsolete
	// brp_commit_wp_response = 3622 // obsolete
	// brp_process_wp_reports = 3623 // obsolete
	// brp_process_payment_rules = 3624 // obsolete
	// brp_process_partner_payments = 3625 // obsolete
	// brp_check_settlement_reports = 3626 // obsolete
	// brp_post_tax_to_avalara = 3628 // obsolete
	brp_post_transaction_tax = 3629
	brp_post_transaction_tax_response = 3630
	// brp_process_im_reports = 3631 // obsolete

	// base_am_range2 = 4000
	am_create_chat = 4001
	am_create_chat_response = 4002
	// am_update_chat_metadata = 4003 // removed
	// am_publish_chat_metadata = 4004 // removed
	am_set_profile_url = 4005
	am_get_account_email_address = 4006
	am_get_account_email_address_response = 4007
	// am_request_friend_data = 4008 // removed "renamed to AMRequestClanData"
	am_request_clan_data = 4008
	am_route_to_clients = 4009
	am_leave_clan = 4010
	am_clan_permissions = 4011
	am_clan_permissions_response = 4012
	// am_create_clan_event = 4013 // obsolete "renamed to AMCreateClanEventDummyForRateLimiting"
	am_create_clan_event_dummy_for_rate_limiting = 4013
	// am_create_clan_event_response = 4014 // obsolete
	// am_update_clan_event = 4015 // obsolete "renamed to AMUpdateClanEventDummyForRateLimiting"
	am_update_clan_event_dummy_for_rate_limiting = 4015
	// am_update_clan_event_response = 4016 // obsolete
	// am_get_clan_events = 4017 // obsolete
	// am_get_clan_events_response = 4018 // obsolete
	// am_delete_clan_event = 4019 // obsolete
	// am_delete_clan_event_response = 4020 // obsolete
	am_set_clan_permission_settings = 4021
	am_set_clan_permission_settings_response = 4022
	am_get_clan_permission_settings = 4023
	am_get_clan_permission_settings_response = 4024
	am_publish_chat_room_info = 4025
	client_chat_room_info = 4026
	// am_create_clan_announcement = 4027 // removed
	// am_create_clan_announcement_response = 4028 // removed
	// am_update_clan_announcement = 4029 // removed
	// am_update_clan_announcement_response = 4030 // removed
	// am_get_clan_announcements_count = 4031 // removed
	// am_get_clan_announcements_count_response = 4032 // removed
	// am_get_clan_announcements = 4033 // removed
	// am_get_clan_announcements_response = 4034 // removed
	// am_delete_clan_announcement = 4035 // removed
	// am_delete_clan_announcement_response = 4036 // removed
	// am_get_single_clan_announcement = 4037 // removed
	// am_get_single_clan_announcement_response = 4038 // removed
	am_get_clan_history = 4039
	am_get_clan_history_response = 4040
	am_get_clan_permission_bits = 4041
	am_get_clan_permission_bits_response = 4042
	am_set_clan_permission_bits = 4043
	am_set_clan_permission_bits_response = 4044
	am_session_info_request = 4045
	am_session_info_response = 4046
	am_validate_wg_token = 4047
	// am_get_single_clan_event = 4048 // obsolete
	// am_get_single_clan_event_response = 4049 // obsolete
	am_get_clan_rank = 4050
	am_get_clan_rank_response = 4051
	am_set_clan_rank = 4052
	am_set_clan_rank_response = 4053
	am_get_clan_potw = 4054
	am_get_clan_potw_response = 4055
	am_set_clan_potw = 4056
	am_set_clan_potw_response = 4057
	// am_request_chat_metadata = 4058 // removed
	am_dump_user = 4059
	am_kick_user_from_clan = 4060
	am_add_founder_to_clan = 4061
	am_validate_wg_token_response = 4062
	// am_set_community_state = 4063 // obsolete
	am_set_account_details = 4064
	am_get_chat_ban_list = 4065
	am_get_chat_ban_list_response = 4066
	am_un_ban_from_chat = 4067
	am_set_clan_details = 4068
	am_get_account_links = 4069
	am_get_account_links_response = 4070
	am_set_account_links = 4071
	am_set_account_links_response = 4072
	// am_get_user_game_stats = 4073 // obsolete "renamed to UGSGetUserGameStats"
	ugs_get_user_game_stats = 4073
	// am_get_user_game_stats_response = 4074 // obsolete "renamed to UGSGetUserGameStatsResponse"
	ugs_get_user_game_stats_response = 4074
	am_check_clan_membership = 4075
	am_get_clan_members = 4076
	am_get_clan_members_response = 4077
	// am_join_public_clan = 4078 // obsolete
	am_notify_chat_of_clan_change = 4079
	am_resubmit_purchase = 4080
	am_add_friend = 4081
	am_add_friend_response = 4082
	am_remove_friend = 4083
	am_dump_clan = 4084
	am_change_clan_owner = 4085
	am_cancel_easy_collect = 4086
	am_cancel_easy_collect_response = 4087
	// am_get_clan_membership_list = 4088 // removed
	// am_get_clan_membership_list_response = 4089 // removed
	am_clans_in_common = 4090
	am_clans_in_common_response = 4091
	am_is_valid_account_id = 4092
	// am_convert_clan = 4093 // obsolete
	// am_get_gift_target_list_relay = 4094 // removed
	am_wipe_friends_list = 4095
	am_set_ignored = 4096
	am_clans_in_common_count_response = 4097
	am_friends_list = 4098
	am_friends_list_response = 4099
	am_friends_in_common = 4100
	am_friends_in_common_response = 4101
	am_friends_in_common_count_response = 4102
	am_clans_in_common_count = 4103
	am_challenge_verdict = 4104
	am_challenge_notification = 4105
	am_find_gs_by_ip = 4106
	am_found_gs_by_ip = 4107
	am_gift_revoked = 4108
	// am_create_account_record = 4109 // obsolete
	am_user_clan_list = 4110
	am_user_clan_list_response = 4111
	am_get_account_details2 = 4112
	am_get_account_details_response2 = 4113
	am_set_community_profile_settings = 4114
	am_set_community_profile_settings_response = 4115
	am_get_community_privacy_state = 4116
	am_get_community_privacy_state_response = 4117
	am_check_clan_invite_rate_limiting = 4118
	// am_get_user_achievement_status = 4119 // obsolete "renamed to UGSGetUserAchievementStatus"
	ugs_get_user_achievement_status = 4119
	am_get_ignored = 4120
	am_get_ignored_response = 4121
	am_set_ignored_response = 4122
	am_set_friend_relationship_none = 4123
	am_get_friend_relationship = 4124
	am_get_friend_relationship_response = 4125
	am_service_modules_cache = 4126
	am_service_modules_call = 4127
	am_service_modules_call_response = 4128
	// am_get_captcha_data_for_ip = 4129 // obsolete
	// am_get_captcha_data_for_ip_response = 4130 // obsolete
	// am_validate_captcha_data_for_ip = 4131 // obsolete
	// am_validate_captcha_data_for_ip_response = 4132 // obsolete
	// am_track_failed_auth_by_ip = 4133 // obsolete
	// am_get_captcha_data_by_gid = 4134 // obsolete
	// am_get_captcha_data_by_gid_response = 4135 // obsolete
	// am_get_lobby_list = 4136 // removed
	// am_get_lobby_list_response = 4137 // removed
	// am_get_lobby_metadata = 4138 // removed
	// am_get_lobby_metadata_response = 4139 // removed
	community_add_friend_news = 4140
	// am_add_clan_news = 4141 // removed
	// am_write_news = 4142 // removed
	am_find_clan_user = 4143
	am_find_clan_user_response = 4144
	am_ban_from_chat = 4145
	// am_get_user_history_response = 4146 // removed
	am_get_user_news_subscriptions = 4147
	am_get_user_news_subscriptions_response = 4148
	am_set_user_news_subscriptions = 4149
	// am_get_user_news = 4150 // removed
	// am_get_user_news_response = 4151 // removed
	am_send_queued_emails = 4152
	am_set_license_flags = 4153
	// am_get_user_history = 4154 // removed
	community_delete_user_news = 4155
	am_allow_user_files_request = 4156
	am_allow_user_files_response = 4157
	am_get_account_status = 4158
	am_get_account_status_response = 4159
	am_edit_ban_reason = 4160
	am_check_clan_membership_response = 4161
	am_probe_clan_membership_list = 4162
	am_probe_clan_membership_list_response = 4163
	ugs_get_user_achievement_status_response = 4164
	am_get_friends_lobbies = 4165
	am_get_friends_lobbies_response = 4166
	am_get_user_friend_news_response = 4172
	community_get_user_friend_news = 4173
	am_get_user_clans_news_response = 4174
	am_get_user_clans_news = 4175
	// am_store_init_purchase = 4176 // removed
	// am_store_init_purchase_response = 4177 // removed
	// am_store_get_final_price = 4178 // removed
	// am_store_get_final_price_response = 4179 // removed
	// am_store_complete_purchase = 4180 // removed
	// am_store_cancel_purchase = 4181 // removed
	// am_store_purchase_response = 4182 // removed
	// am_create_account_record_in_steam3 = 4183 // removed
	am_get_previous_cb_account = 4184
	am_get_previous_cb_account_response = 4185
	// am_update_billing_address = 4186 // removed
	// am_update_billing_address_response = 4187 // removed
	// am_get_billing_address = 4188 // removed
	// am_get_billing_address_response = 4189 // removed
	am_get_user_license_history = 4190
	am_get_user_license_history_response = 4191
	am_support_change_password = 4194
	am_support_change_email = 4195
	// am_support_change_secret_qa = 4196 // removed
	am_reset_user_verification_gs_by_ip = 4197
	am_update_gs_play_stats = 4198
	am_support_enable_or_disable = 4199
	// am_get_comments = 4200 // removed
	// am_get_comments_response = 4201 // removed
	// am_add_comment = 4202 // removed
	// am_add_comment_response = 4203 // removed
	// am_delete_comment = 4204 // removed
	// am_delete_comment_response = 4205 // removed
	am_get_purchase_status = 4206
	am_support_is_account_enabled = 4209
	am_support_is_account_enabled_response = 4210
	// am_get_user_stats = 4211 // obsolete "renamed to UGSGetUserStats"
	ugs_get_user_stats = 4211
	am_support_kick_session = 4212
	amgs_search = 4213
	marketing_message_update = 4216
	// am_route_friend_msg = 4219 // obsolete "renamed to ChatServerRouteFriendMsg"
	chat_server_route_friend_msg = 4219
	am_ticket_auth_request_or_response = 4220
	am_verify_depot_management_rights = 4222
	am_verify_depot_management_rights_response = 4223
	am_add_free_license = 4224
	// am_get_user_friends_minutes_played = 4225 // removed
	// am_get_user_friends_minutes_played_response = 4226 // removed
	// am_get_user_minutes_played = 4227 // removed
	// am_get_user_minutes_played_response = 4228 // removed
	am_validate_email_link = 4231
	am_validate_email_link_response = 4232
	// am_add_users_to_marketing_treatment = 4234 // removed
	// am_store_user_stats = 4236 // obsolete "renamed to UGSStoreUserStats"
	ugs_store_user_stats = 4236
	// am_get_user_gameplay_info = 4237 // removed
	// am_get_user_gameplay_info_response = 4238 // removed
	// am_get_card_list = 4239 // removed
	// am_get_card_list_response = 4240 // removed
	am_delete_stored_card = 4241
	am_revoke_legacy_game_keys = 4242
	am_get_wallet_details = 4244
	am_get_wallet_details_response = 4245
	am_delete_stored_payment_info = 4246
	am_get_stored_payment_summary = 4247
	am_get_stored_payment_summary_response = 4248
	am_get_wallet_conversion_rate = 4249
	am_get_wallet_conversion_rate_response = 4250
	am_convert_wallet = 4251
	am_convert_wallet_response = 4252
	// am_relay_get_friends_who_play_game = 4253 // removed
	// am_relay_get_friends_who_play_game_response = 4254 // removed
	am_set_pre_approval = 4255
	am_set_pre_approval_response = 4256
	// am_marketing_treatment_update = 4257 // removed
	am_create_refund = 4258
	// am_create_refund_response = 4259 // obsolete
	am_create_chargeback = 4260
	// am_create_chargeback_response = 4261 // obsolete
	am_create_dispute = 4262
	// am_create_dispute_response = 4263 // obsolete
	am_clear_dispute = 4264
	// am_clear_dispute_response = 4265 // obsolete "renamed to AMCreateFinancialAdjustment"
	am_create_financial_adjustment = 4265
	am_player_nickname_list = 4266
	am_player_nickname_list_response = 4267
	am_set_drm_test_config = 4268
	am_get_user_current_game_info = 4269
	am_get_user_current_game_info_response = 4270
	am_get_gs_player_list = 4271
	am_get_gs_player_list_response = 4272
	// am_update_persona_state_cache = 4275 // removed
	am_get_game_members = 4276
	am_get_game_members_response = 4277
	am_get_steam_id_for_micro_txn = 4278
	am_get_steam_id_for_micro_txn_response = 4279
	// am_add_publisher_user = 4280 // obsolete "renamed to AMSetPartnerMember"
	am_set_partner_member = 4280
	am_remove_publisher_user = 4281
	am_get_user_license_list = 4282
	am_get_user_license_list_response = 4283
	am_reload_game_group_policy = 4284
	am_add_free_license_response = 4285
	amvac_status_update = 4286
	am_get_account_details = 4287
	am_get_account_details_response = 4288
	am_get_player_link_details = 4289
	am_get_player_link_details_response = 4290
	// am_subscribe_to_persona_feed = 4291 // removed
	// am_get_user_vac_ban_list = 4292 // removed
	// am_get_user_vac_ban_list_response = 4293 // removed
	am_get_account_flags_for_wg_spoofing = 4294
	am_get_account_flags_for_wg_spoofing_response = 4295
	// am_get_friends_wishlist_info = 4296 // removed
	// am_get_friends_wishlist_info_response = 4297 // removed
	am_get_clan_officers = 4298
	am_get_clan_officers_response = 4299
	am_name_change = 4300
	am_get_name_history = 4301
	am_get_name_history_response = 4302
	am_update_provider_status = 4305
	// am_clear_persona_metadata_blob = 4306 // removed
	am_support_remove_account_security = 4307
	am_is_account_in_captcha_grace_period = 4308
	am_is_account_in_captcha_grace_period_response = 4309
	am_account_ps3_unlink = 4310
	am_account_ps3_unlink_response = 4311
	// am_store_user_stats_response = 4312 // obsolete "renamed to UGSStoreUserStatsResponse"
	ugs_store_user_stats_response = 4312
	am_get_account_psn_info = 4313
	am_get_account_psn_info_response = 4314
	am_authenticated_player_list = 4315
	am_get_user_gifts = 4316
	am_get_user_gifts_response = 4317
	am_transfer_locked_gifts = 4320
	am_transfer_locked_gifts_response = 4321
	am_player_hosted_on_game_server = 4322
	am_get_account_ban_info = 4323
	am_get_account_ban_info_response = 4324
	am_record_ban_enforcement = 4325
	am_rollback_gift_transfer = 4326
	am_rollback_gift_transfer_response = 4327
	am_handle_pending_transaction = 4328
	am_request_clan_details = 4329
	am_delete_stored_paypal_agreement = 4330
	am_game_server_update = 4331
	am_game_server_remove = 4332
	am_get_paypal_agreements = 4333
	am_get_paypal_agreements_response = 4334
	am_game_server_player_compatibility_check = 4335
	am_game_server_player_compatibility_check_response = 4336
	am_renew_license = 4337
	am_get_account_community_ban_info = 4338
	am_get_account_community_ban_info_response = 4339
	am_game_server_account_change_password = 4340
	am_game_server_account_delete_account = 4341
	am_renew_agreement = 4342
	// am_send_email = 4343 // removed
	am_xsolla_payment = 4344
	am_xsolla_payment_response = 4345
	am_acct_allowed_to_purchase = 4346
	am_acct_allowed_to_purchase_response = 4347
	am_swap_kiosk_deposit = 4348
	am_swap_kiosk_deposit_response = 4349
	am_set_user_gift_unowned = 4350
	am_set_user_gift_unowned_response = 4351
	am_claim_unowned_user_gift = 4352
	am_claim_unowned_user_gift_response = 4353
	am_set_clan_name = 4354
	am_set_clan_name_response = 4355
	am_grant_coupon = 4356
	am_grant_coupon_response = 4357
	am_is_package_restricted_in_user_country = 4358
	am_is_package_restricted_in_user_country_response = 4359
	am_handle_pending_transaction_response = 4360
	am_grant_guest_passes2 = 4361
	am_grant_guest_passes2_response = 4362
	// am_session_query = 4363 // obsolete
	// am_session_query_response = 4364 // obsolete
	am_get_player_ban_details = 4365
	am_get_player_ban_details_response = 4366
	am_finalize_purchase = 4367
	am_finalize_purchase_response = 4368
	am_persona_change_response = 4372
	am_get_clan_details_for_forum_creation = 4373
	am_get_clan_details_for_forum_creation_response = 4374
	am_get_pending_notification_count = 4375
	am_get_pending_notification_count_response = 4376
	am_password_hash_upgrade = 4377
	// am_mo_pay_payment = 4378 // obsolete
	// am_mo_pay_payment_response = 4379 // obsolete
	am_boa_compra_payment = 4380
	am_boa_compra_payment_response = 4381
	// am_expire_captcha_by_gid = 4382 // obsolete
	am_complete_external_purchase = 4383
	am_complete_external_purchase_response = 4384
	am_resolve_negative_wallet_credits = 4385
	am_resolve_negative_wallet_credits_response = 4386
	// am_payelp_payment = 4387 // obsolete
	// am_payelp_payment_response = 4388 // obsolete
	am_player_get_clan_basic_details = 4389
	am_player_get_clan_basic_details_response = 4390
	ammol_payment = 4391
	ammol_payment_response = 4392
	get_user_ip_country = 4393
	get_user_ip_country_response = 4394
	notification_of_suspicious_activity = 4395
	am_degica_payment = 4396
	am_degica_payment_response = 4397
	ame_club_payment = 4398
	ame_club_payment_response = 4399
	am_pay_pal_payments_hub_payment = 4400
	am_pay_pal_payments_hub_payment_response = 4401
	am_two_factor_recover_authenticator_request = 4402
	am_two_factor_recover_authenticator_response = 4403
	am_smart2_pay_payment = 4404
	am_smart2_pay_payment_response = 4405
	am_validate_password_reset_code_and_send_sms_request = 4406
	am_validate_password_reset_code_and_send_sms_response = 4407
	am_get_account_reset_details_request = 4408
	am_get_account_reset_details_response = 4409
	am_bit_pay_payment = 4410
	am_bit_pay_payment_response = 4411
	am_send_account_info_update = 4412
	am_send_scheduled_gift = 4413
	am_nodwin_payment = 4414
	am_nodwin_payment_response = 4415
	am_resolve_wallet_revoke = 4416
	am_resolve_wallet_reverse_revoke = 4417
	am_funded_payment = 4418
	am_funded_payment_response = 4419
	am_request_persona_update_for_chat_server = 4420
	am_perfect_world_payment = 4421
	am_perfect_world_payment_response = 4422

	// base_ps_range = 5000
	ps_create_shopping_cart = 5001
	ps_create_shopping_cart_response = 5002
	ps_is_valid_shopping_cart = 5003
	ps_is_valid_shopping_cart_response = 5004
	ps_add_package_to_shopping_cart = 5005
	ps_add_package_to_shopping_cart_response = 5006
	ps_remove_line_item_from_shopping_cart = 5007
	ps_remove_line_item_from_shopping_cart_response = 5008
	ps_get_shopping_cart_contents = 5009
	ps_get_shopping_cart_contents_response = 5010
	ps_add_wallet_credit_to_shopping_cart = 5011
	ps_add_wallet_credit_to_shopping_cart_response = 5012

	// base_ufs_range = 5200
	client_ufs_upload_file_request = 5202
	client_ufs_upload_file_response = 5203
	client_ufs_upload_file_chunk = 5204
	client_ufs_upload_file_finished = 5205
	client_ufs_get_file_list_for_app = 5206
	client_ufs_get_file_list_for_app_response = 5207
	client_ufs_download_request = 5210
	client_ufs_download_response = 5211
	client_ufs_download_chunk = 5212
	client_ufs_login_request = 5213
	client_ufs_login_response = 5214
	ufs_reload_partition_info = 5215
	client_ufs_transfer_heartbeat = 5216
	ufs_synchronize_file = 5217
	ufs_synchronize_file_response = 5218
	client_ufs_delete_file_request = 5219
	client_ufs_delete_file_response = 5220
	// ufs_download_request = 5221 // removed
	// ufs_download_response = 5222 // removed
	// ufs_download_chunk = 5223 // removed
	client_ufs_get_ugc_details = 5226
	client_ufs_get_ugc_details_response = 5227
	ufs_update_file_flags = 5228
	ufs_update_file_flags_response = 5229
	client_ufs_get_single_file_info = 5230
	client_ufs_get_single_file_info_response = 5231
	client_ufs_share_file = 5232
	client_ufs_share_file_response = 5233
	ufs_reload_account = 5234
	ufs_reload_account_response = 5235
	ufs_update_record_batched = 5236
	ufs_update_record_batched_response = 5237
	ufs_migrate_file = 5238
	ufs_migrate_file_response = 5239
	ufs_get_ugcur_ls = 5240
	ufs_get_ugcur_ls_response = 5241
	ufs_http_upload_file_finish_request = 5242
	ufs_http_upload_file_finish_response = 5243
	ufs_download_start_request = 5244
	ufs_download_start_response = 5245
	ufs_download_chunk_request = 5246
	ufs_download_chunk_response = 5247
	ufs_download_finish_request = 5248
	ufs_download_finish_response = 5249
	ufs_flush_url_cache = 5250
	// ufs_upload_commit = 5251 // obsolete "renamed to ClientUFSUploadCommit"
	client_ufs_upload_commit = 5251
	// ufs_upload_commit_response = 5252 // obsolete "renamed to ClientUFSUploadCommitResponse"
	client_ufs_upload_commit_response = 5252
	ufs_migrate_file_app_id = 5253
	ufs_migrate_file_app_id_response = 5254

	// base_client2 = 5400
	client_request_forgotten_password_email = 5401
	client_request_forgotten_password_email_response = 5402
	client_create_account_response = 5403
	client_reset_forgotten_password = 5404
	client_reset_forgotten_password_response = 5405
	// client_create_account2 = 5406 // obsolete
	client_inform_of_reset_forgotten_password = 5407
	client_inform_of_reset_forgotten_password_response = 5408
	// client_anon_user_log_on_deprecated = 5409 // removed
	client_games_played_with_data_blob = 5410
	client_update_user_game_info = 5411
	client_file_to_download = 5412
	client_file_to_download_response = 5413
	client_lbs_set_score = 5414
	client_lbs_set_score_response = 5415
	client_lbs_find_or_create_lb = 5416
	client_lbs_find_or_create_lb_response = 5417
	client_lbs_get_lb_entries = 5418
	client_lbs_get_lb_entries_response = 5419
	// client_marketing_message_update = 5420 // removed
	client_chat_declined = 5426
	client_friend_msg_incoming = 5427
	// client_auth_list_deprecated = 5428 // removed
	client_ticket_auth_complete = 5429
	client_is_limited_account = 5430
	client_request_auth_list = 5431
	client_auth_list = 5432
	client_stat = 5433
	client_p2_p_connection_info = 5434
	client_p2_p_connection_fail_info = 5435
	// client_get_number_of_current_players = 5436 // removed
	// client_get_number_of_current_players_response = 5437 // removed
	client_get_depot_decryption_key = 5438
	client_get_depot_decryption_key_response = 5439
	gs_perform_hardware_survey = 5440
	// client_get_app_beta_passwords = 5441 // removed
	// client_get_app_beta_passwords_response = 5442 // removed
	client_enable_test_license = 5443
	client_enable_test_license_response = 5444
	client_disable_test_license = 5445
	client_disable_test_license_response = 5446
	client_request_validation_mail = 5448
	client_request_validation_mail_response = 5449
	client_check_app_beta_password = 5450
	client_check_app_beta_password_response = 5451
	client_to_gc = 5452
	client_from_gc = 5453
	client_request_change_mail = 5454
	client_request_change_mail_response = 5455
	client_email_addr_info = 5456
	client_password_change3 = 5457
	client_email_change3 = 5458
	client_personal_qa_change3 = 5459
	client_reset_forgotten_password3 = 5460
	client_request_forgotten_password_email3 = 5461
	// client_create_account3 = 5462 // removed
	client_new_login_key = 5463
	client_new_login_key_accepted = 5464
	// client_log_on_with_hash_deprecated = 5465 // removed
	client_store_user_stats2 = 5466
	client_stats_updated = 5467
	client_activate_oem_license = 5468
	client_register_oem_machine = 5469
	client_register_oem_machine_response = 5470
	client_requested_client_stats = 5480
	client_stat2_int32 = 5481
	client_stat2 = 5482
	client_verify_password = 5483
	client_verify_password_response = 5484
	client_drm_download_request = 5485
	client_drm_download_response = 5486
	client_drm_final_result = 5487
	client_get_friends_who_play_game = 5488
	client_get_friends_who_play_game_response = 5489
	client_ogs_begin_session = 5490
	client_ogs_begin_session_response = 5491
	client_ogs_end_session = 5492
	client_ogs_end_session_response = 5493
	client_ogs_write_row = 5494
	client_drm_test = 5495
	client_drm_test_result = 5496
	client_server_unavailable = 5500
	client_servers_available = 5501
	client_register_auth_ticket_with_cm = 5502
	client_gc_msg_failed = 5503
	client_micro_txn_auth_request = 5504
	client_micro_txn_authorize = 5505
	client_micro_txn_authorize_response = 5506
	client_app_minutes_played_data = 5507
	client_get_micro_txn_info = 5508
	client_get_micro_txn_info_response = 5509
	client_marketing_message_update2 = 5510
	client_deregister_with_server = 5511
	client_subscribe_to_persona_feed = 5512
	client_logon = 5514
	client_get_client_details = 5515
	client_get_client_details_response = 5516
	client_report_overlay_detour_failure = 5517
	client_get_client_app_list = 5518
	client_get_client_app_list_response = 5519
	client_install_client_app = 5520
	client_install_client_app_response = 5521
	client_uninstall_client_app = 5522
	client_uninstall_client_app_response = 5523
	client_set_client_app_update_state = 5524
	client_set_client_app_update_state_response = 5525
	client_request_encrypted_app_ticket = 5526
	client_request_encrypted_app_ticket_response = 5527
	client_wallet_info_update = 5528
	client_lbs_set_ugc = 5529
	client_lbs_set_ugc_response = 5530
	client_am_get_clan_officers = 5531
	client_am_get_clan_officers_response = 5532
	// client_check_file_signature = 5533 // removed
	// client_check_file_signature_response = 5534 // removed
	client_friend_profile_info = 5535
	client_friend_profile_info_response = 5536
	client_update_machine_auth = 5537
	client_update_machine_auth_response = 5538
	client_read_machine_auth = 5539
	client_read_machine_auth_response = 5540
	client_request_machine_auth = 5541
	client_request_machine_auth_response = 5542
	client_screenshots_changed = 5543
	// client_email_change4 = 5544 // obsolete
	// client_email_change_response4 = 5545 // obsolete
	client_get_cdn_auth_token = 5546
	client_get_cdn_auth_token_response = 5547
	client_download_rate_statistics = 5548
	client_request_account_data = 5549
	client_request_account_data_response = 5550
	client_reset_forgotten_password4 = 5551
	client_hide_friend = 5552
	client_friends_groups_list = 5553
	client_get_clan_activity_counts = 5554
	client_get_clan_activity_counts_response = 5555
	client_ogs_report_string = 5556
	client_ogs_report_bug = 5557
	client_sent_logs = 5558
	client_logon_game_server = 5559
	am_client_create_friends_group = 5560
	am_client_create_friends_group_response = 5561
	am_client_delete_friends_group = 5562
	am_client_delete_friends_group_response = 5563
	// am_client_rename_friends_group = 5564 // obsolete "renamed to AMClientManageFriendsGroup"
	am_client_manage_friends_group = 5564
	// am_client_rename_friends_group_response = 5565 // obsolete "renamed to AMClientManageFriendsGroupResponse"
	am_client_manage_friends_group_response = 5565
	am_client_add_friend_to_group = 5566
	am_client_add_friend_to_group_response = 5567
	am_client_remove_friend_from_group = 5568
	am_client_remove_friend_from_group_response = 5569
	client_am_get_persona_name_history = 5570
	client_am_get_persona_name_history_response = 5571
	client_request_free_license = 5572
	client_request_free_license_response = 5573
	client_drm_download_request_with_crash_data = 5574
	client_auth_list_ack = 5575
	client_item_announcements = 5576
	client_request_item_announcements = 5577
	client_friend_msg_echo_to_sender = 5578
	// client_change_steam_guard_options = 5579 // removed
	// client_change_steam_guard_options_response = 5580 // removed
	client_ogs_game_server_ping_sample = 5581
	client_comment_notifications = 5582
	client_request_comment_notifications = 5583
	client_persona_change_response = 5584
	client_request_web_api_authenticate_user_nonce = 5585
	client_request_web_api_authenticate_user_nonce_response = 5586
	client_player_nickname_list = 5587
	am_client_set_player_nickname = 5588
	am_client_set_player_nickname_response = 5589
	// client_request_o_auth_token_for_app = 5590 // removed
	// client_request_o_auth_token_for_app_response = 5591 // removed
	// client_create_account_proto = 5590 // obsolete
	// client_create_account_proto_response = 5591 // obsolete
	client_get_number_of_current_players_dp = 5592
	client_get_number_of_current_players_dp_response = 5593
	// client_service_method = 5594 // obsolete "renamed to ClientServiceMethodLegacy"
	client_service_method_legacy = 5594
	// client_service_method_response = 5595 // obsolete "renamed to ClientServiceMethodLegacyResponse"
	client_service_method_legacy_response = 5595
	client_friend_user_status_published = 5596
	client_current_ui_mode = 5597
	client_vanity_url_changed_notification = 5598
	client_user_notifications = 5599

	// base_dfs = 5600
	dfs_get_file = 5601
	dfs_install_local_file = 5602
	dfs_connection = 5603
	dfs_connection_reply = 5604
	client_dfs_authenticate_request = 5605
	client_dfs_authenticate_response = 5606
	client_dfs_end_session = 5607
	dfs_purge_file = 5608
	dfs_route_file = 5609
	dfs_get_file_from_server = 5610
	dfs_accepted_response = 5611
	dfs_request_pingback = 5612
	dfs_recv_transmit_file = 5613
	dfs_send_transmit_file = 5614
	dfs_request_pingback2 = 5615
	dfs_response_pingback2 = 5616
	client_dfs_download_status = 5617
	dfs_start_transfer = 5618
	dfs_transfer_complete = 5619
	dfs_route_file_response = 5620
	client_networking_cert_request = 5621
	client_networking_cert_request_response = 5622
	client_challenge_request = 5623
	client_challenge_response = 5624
	badge_crafted_notification = 5625
	client_networking_mobile_cert_request = 5626
	client_networking_mobile_cert_request_response = 5627

	// base_mds = 5800
	// client_mds_login_request = 5801 // removed
	// client_mds_login_response = 5802 // removed
	// client_mds_upload_manifest_request = 5803 // removed
	// client_mds_upload_manifest_response = 5804 // removed
	// client_mds_transmit_manifest_data_chunk = 5805 // removed
	// client_mds_heartbeat = 5806 // removed
	// client_mds_upload_depot_chunks = 5807 // removed
	// client_mds_upload_depot_chunks_response = 5808 // removed
	// client_mds_init_depot_build_request = 5809 // removed
	// client_mds_init_depot_build_response = 5810 // removed
	am_to_mds_get_depot_decryption_key = 5812
	mds_to_am_get_depot_decryption_key_response = 5813
	// mds_get_versions_for_depot = 5814 // removed
	// mds_get_versions_for_depot_response = 5815 // removed
	// mds_set_public_version_for_depot = 5816 // removed
	// mds_set_public_version_for_depot_response = 5817 // removed
	// client_mds_init_workshop_build_request = 5816 // removed
	// client_mds_init_workshop_build_response = 5817 // removed
	// client_mds_get_depot_manifest = 5818 // removed
	// client_mds_get_depot_manifest_response = 5819 // removed
	// client_mds_get_depot_manifest_chunk = 5820 // removed
	// client_mds_upload_rate_test = 5823 // removed
	// client_mds_upload_rate_test_response = 5824 // removed
	// mds_download_depot_chunks_ack = 5825 // removed
	// mds_content_server_stats_broadcast = 5826 // removed
	mds_content_server_config_request = 5827
	mds_content_server_config = 5828
	mds_get_depot_manifest = 5829
	mds_get_depot_manifest_response = 5830
	mds_get_depot_manifest_chunk = 5831
	mds_get_depot_chunk = 5832
	mds_get_depot_chunk_response = 5833
	mds_get_depot_chunk_chunk = 5834
	// mds_update_content_server_config = 5835 // removed
	// mds_get_server_list_for_user = 5836 // obsolete
	// mds_get_server_list_for_user_response = 5837 // obsolete
	// client_mds_register_app_build = 5838 // removed
	// client_mds_register_app_build_response = 5839 // removed
	// client_mds_set_app_build_live = 5840 // removed
	// client_mds_set_app_build_live_response = 5841 // removed
	// client_mds_get_prev_depot_build = 5842 // removed
	// client_mds_get_prev_depot_build_response = 5843 // removed
	mds_to_cs_flush_chunk = 5844
	// client_mds_sign_install_script = 5845 // removed
	// client_mds_sign_install_script_response = 5846 // removed
	mds_migrate_chunk = 5847
	mds_migrate_chunk_response = 5848
	mds_to_cs_flush_manifest = 5849

	// cs_base = 6200
	cs_ping = 6201
	cs_ping_response = 6202

	// gms_base = 6400
	gms_game_server_replicate = 6401
	client_gms_server_query = 6403
	gms_client_server_query_response = 6404
	amgms_game_server_update = 6405
	amgms_game_server_remove = 6406
	game_server_out_of_date = 6407

	// device_authorization_base = 6500
	client_authorize_local_device_request = 6501
	// client_authorize_local_device = 6502 // removed
	client_authorize_local_device_response = 6502
	client_deauthorize_device_request = 6503
	client_deauthorize_device = 6504
	client_use_local_device_authorizations = 6505
	client_get_authorized_devices = 6506
	client_get_authorized_devices_response = 6507
	am_notify_session_device_authorized = 6508
	client_authorize_local_device_notification = 6509

	// mms_base = 6600
	client_mms_create_lobby = 6601
	client_mms_create_lobby_response = 6602
	client_mms_join_lobby = 6603
	client_mms_join_lobby_response = 6604
	client_mms_leave_lobby = 6605
	client_mms_leave_lobby_response = 6606
	client_mms_get_lobby_list = 6607
	client_mms_get_lobby_list_response = 6608
	client_mms_set_lobby_data = 6609
	client_mms_set_lobby_data_response = 6610
	client_mms_get_lobby_data = 6611
	client_mms_lobby_data = 6612
	client_mms_send_lobby_chat_msg = 6613
	client_mms_lobby_chat_msg = 6614
	client_mms_set_lobby_owner = 6615
	client_mms_set_lobby_owner_response = 6616
	client_mms_set_lobby_game_server = 6617
	client_mms_lobby_game_server_set = 6618
	client_mms_user_joined_lobby = 6619
	client_mms_user_left_lobby = 6620
	client_mms_invite_to_lobby = 6621
	client_mms_flush_frenemy_list_cache = 6622
	client_mms_flush_frenemy_list_cache_response = 6623
	client_mms_set_lobby_linked = 6624
	client_mms_set_ratelimit_policy_on_client = 6625
	client_mms_get_lobby_status = 6626
	client_mms_get_lobby_status_response = 6627
	mms_get_lobby_list = 6628
	mms_get_lobby_list_response = 6629

	// non_std_msg_base = 6800
	non_std_msg_memcached = 6801
	non_std_msg_http_server = 6802
	non_std_msg_http_client = 6803
	non_std_msg_wg_response = 6804
	non_std_msg_php_simulator = 6805
	non_std_msg_chase = 6806
	non_std_msg_dfs_transfer = 6807
	non_std_msg_tests = 6808
	non_std_msg_um_qpipe_aapl = 6809
	non_std_msg_syslog = 6810
	non_std_msg_logsink = 6811
	non_std_msg_steam2_emulator = 6812
	non_std_msg_rtmp_server = 6813
	non_std_msg_web_socket = 6814
	non_std_msg_redis = 6815

	// uds_base = 7000
	client_udsp2_p_session_started = 7001
	client_udsp2_p_session_ended = 7002
	uds_render_user_auth = 7003
	uds_render_user_auth_response = 7004
	// client_uds_invite_to_game = 7005 // obsolete "renamed to ClientInviteToGame"
	client_invite_to_game = 7005
	// uds_find_session = 7006 // removed "renamed to UDSHasSession"
	uds_has_session = 7006
	// uds_find_session_response = 7007 // removed "renamed to UDSHasSessionResponse"
	uds_has_session_response = 7007

	// mpas_base = 7100
	mpas_vac_ban_reset = 7101

	// kgs_base = 7200
	// kgs_allocate_key_range = 7201 // removed
	// kgs_allocate_key_range_response = 7202 // removed
	// kgs_generate_keys = 7203 // removed
	// kgs_generate_keys_response = 7204 // removed
	// kgs_remap_keys = 7205 // removed
	// kgs_remap_keys_response = 7206 // removed
	// kgs_generate_game_stop_wc_keys = 7207 // removed
	// kgs_generate_game_stop_wc_keys_response = 7208 // removed

	// ucm_base = 7300
	client_ucm_add_screenshot = 7301
	client_ucm_add_screenshot_response = 7302
	// ucm_validate_object_exists = 7303 // removed
	// ucm_validate_object_exists_response = 7304 // removed
	ucm_reset_community_content = 7307
	ucm_reset_community_content_response = 7308
	client_ucm_delete_screenshot = 7309
	client_ucm_delete_screenshot_response = 7310
	client_ucm_publish_file = 7311
	client_ucm_publish_file_response = 7312
	// client_ucm_get_published_file_details = 7313 // removed
	// client_ucm_get_published_file_details_response = 7314 // removed
	client_ucm_delete_published_file = 7315
	client_ucm_delete_published_file_response = 7316
	client_ucm_enumerate_user_published_files = 7317
	client_ucm_enumerate_user_published_files_response = 7318
	// client_ucm_subscribe_published_file = 7319 // removed
	// client_ucm_subscribe_published_file_response = 7320 // removed
	client_ucm_enumerate_user_subscribed_files = 7321
	client_ucm_enumerate_user_subscribed_files_response = 7322
	// client_ucm_unsubscribe_published_file = 7323 // removed
	// client_ucm_unsubscribe_published_file_response = 7324 // removed
	client_ucm_update_published_file = 7325
	client_ucm_update_published_file_response = 7326
	ucm_update_published_file = 7327
	ucm_update_published_file_response = 7328
	ucm_delete_published_file = 7329
	ucm_delete_published_file_response = 7330
	ucm_update_published_file_stat = 7331
	// ucm_update_published_file_ban = 7332 // obsolete
	// ucm_update_published_file_ban_response = 7333 // obsolete
	// ucm_update_tagged_screenshot = 7334 // removed
	// ucm_add_tagged_screenshot = 7335 // removed
	// ucm_remove_tagged_screenshot = 7336 // removed
	ucm_reload_published_file = 7337
	ucm_reload_user_file_list_caches = 7338
	ucm_published_file_reported = 7339
	// ucm_update_published_file_incompatible_status = 7340 // obsolete
	ucm_published_file_preview_add = 7341
	ucm_published_file_preview_add_response = 7342
	ucm_published_file_preview_remove = 7343
	ucm_published_file_preview_remove_response = 7344
	// ucm_published_file_preview_change_sort_order = 7345 // removed
	// ucm_published_file_preview_change_sort_order_response = 7346 // removed
	client_ucm_published_file_subscribed = 7347
	client_ucm_published_file_unsubscribed = 7348
	ucm_published_file_subscribed = 7349
	ucm_published_file_unsubscribed = 7350
	ucm_publish_file = 7351
	ucm_publish_file_response = 7352
	ucm_published_file_child_add = 7353
	ucm_published_file_child_add_response = 7354
	ucm_published_file_child_remove = 7355
	ucm_published_file_child_remove_response = 7356
	// ucm_published_file_child_change_sort_order = 7357 // removed
	// ucm_published_file_child_change_sort_order_response = 7358 // removed
	ucm_published_file_parent_changed = 7359
	client_ucm_get_published_files_for_user = 7360
	client_ucm_get_published_files_for_user_response = 7361
	// ucm_get_published_files_for_user = 7362 // removed
	// ucm_get_published_files_for_user_response = 7363 // removed
	client_ucm_set_user_published_file_action = 7364
	client_ucm_set_user_published_file_action_response = 7365
	client_ucm_enumerate_published_files_by_user_action = 7366
	client_ucm_enumerate_published_files_by_user_action_response = 7367
	client_ucm_published_file_deleted = 7368
	ucm_get_user_subscribed_files = 7369
	ucm_get_user_subscribed_files_response = 7370
	ucm_fix_stats_published_file = 7371
	// ucm_delete_old_screenshot = 7372 // removed
	// ucm_delete_old_screenshot_response = 7373 // removed
	// ucm_delete_old_video = 7374 // removed
	// ucm_delete_old_video_response = 7375 // removed
	// ucm_update_old_screenshot_privacy = 7376 // removed
	// ucm_update_old_screenshot_privacy_response = 7377 // removed
	client_ucm_enumerate_user_subscribed_files_with_updates = 7378
	client_ucm_enumerate_user_subscribed_files_with_updates_response = 7379
	ucm_published_file_content_updated = 7380
	// ucm_published_file_updated = 7381 // obsolete "renamed to ClientUCMPublishedFileUpdated"
	client_ucm_published_file_updated = 7381
	client_workshop_item_changes_request = 7382
	client_workshop_item_changes_response = 7383
	client_workshop_item_info_request = 7384
	client_workshop_item_info_response = 7385

	// fs_base = 7500
	client_rich_presence_upload = 7501
	client_rich_presence_request = 7502
	client_rich_presence_info = 7503
	fs_rich_presence_request = 7504
	fs_rich_presence_response = 7505
	fs_compute_frenematrix = 7506
	fs_compute_frenematrix_response = 7507
	fs_play_status_notification = 7508
	// fs_publish_persona_status = 7509 // obsolete
	fs_add_or_remove_follower = 7510
	fs_add_or_remove_follower_response = 7511
	fs_update_following_list = 7512
	fs_comment_notification = 7513
	fs_comment_notification_viewed = 7514
	client_fs_get_follower_count = 7515
	client_fs_get_follower_count_response = 7516
	client_fs_get_is_following = 7517
	client_fs_get_is_following_response = 7518
	client_fs_enumerate_following_list = 7519
	client_fs_enumerate_following_list_response = 7520
	fs_get_pending_notification_count = 7521
	fs_get_pending_notification_count_response = 7522
	// client_fs_offline_message_notification = 7523 // obsolete "Renamed to ClientChatOfflineMessageNotification"
	// client_fs_request_offline_message_count = 7524 // obsolete "Renamed to ClientChatRequestOfflineMessageCount"
	// client_fs_get_friend_message_history = 7525 // obsolete "Renamed to ClientChatGetFriendMessageHistory"
	// client_fs_get_friend_message_history_response = 7526 // obsolete "Renamed to ClientChatGetFriendMessageHistoryResponse"
	// client_fs_get_friend_message_history_for_offline_messages = 7527 // obsolete "Renamed to ClientChatGetFriendMessageHistoryForOfflineMessages"
	client_chat_offline_message_notification = 7523
	client_chat_request_offline_message_count = 7524
	client_chat_get_friend_message_history = 7525
	client_chat_get_friend_message_history_response = 7526
	client_chat_get_friend_message_history_for_offline_messages = 7527
	client_fs_get_friends_steam_levels = 7528
	client_fs_get_friends_steam_levels_response = 7529
	// fs_request_friend_data = 7530 // obsolete "renamed to AMRequestFriendData"
	am_request_friend_data = 7530

	// drm_range2 = 7600
	ceg_version_set_enable_disable_request = 7600
	ceg_version_set_enable_disable_response = 7601
	ceg_prop_status_drms_request = 7602
	ceg_prop_status_drms_response = 7603
	ceg_whack_failure_report_request = 7604
	ceg_whack_failure_report_response = 7605
	drms_fetch_version_set = 7606
	drms_fetch_version_set_response = 7607

	// econ_base = 7700
	econ_trading_initiate_trade_request = 7701
	econ_trading_initiate_trade_proposed = 7702
	econ_trading_initiate_trade_response = 7703
	econ_trading_initiate_trade_result = 7704
	econ_trading_start_session = 7705
	econ_trading_cancel_trade_request = 7706
	econ_flush_inventory_cache = 7707
	econ_flush_inventory_cache_response = 7708
	econ_cd_key_process_transaction = 7711
	econ_cd_key_process_transaction_response = 7712
	econ_get_error_logs = 7713
	econ_get_error_logs_response = 7714

	// rm_range = 7800
	rm_test_verisign_otp = 7800
	rm_test_verisign_otp_response = 7801
	rm_delete_memcached_keys = 7803
	rm_remote_invoke = 7804
	bad_login_ip_list = 7805
	rm_msg_trace_add_trigger = 7806
	rm_msg_trace_remove_trigger = 7807
	rm_msg_trace_event = 7808

	// ugs_base = 7900
	ugs_update_global_stats = 7900
	client_ugs_get_global_stats = 7901
	client_ugs_get_global_stats_response = 7902

	// store_base = 8000
	// store_update_recommendation_count = 8000 // removed

	// umq_base = 8100
	umq_logon_request = 8100
	umq_logon_response = 8101
	umq_logoff_request = 8102
	umq_logoff_response = 8103
	umq_send_chat_message = 8104
	umq_incoming_chat_message = 8105
	umq_poll = 8106
	umq_poll_results = 8107
	umq2_am_client_msg_batch = 8108
	// umq_enqueue_mobile_sale_promotions = 8109 // removed
	// umq_enqueue_mobile_announcements = 8110 // removed

	// workshop_base = 8200
	// workshop_accept_tos_request = 8200 // removed
	// workshop_accept_tos_response = 8201 // removed

	// web_api_base = 8300
	web_api_validate_o_auth2_token = 8300
	web_api_validate_o_auth2_token_response = 8301
	// web_api_invalidate_tokens_for_account = 8302 // removed
	web_api_register_gc_interfaces = 8303
	web_api_invalidate_o_auth_client_cache = 8304
	web_api_invalidate_o_auth_token_cache = 8305
	web_api_set_secrets = 8306

	// backpack_base = 8400
	backpack_add_to_currency = 8401
	backpack_add_to_currency_response = 8402

	// cre_base = 8500
	// cre_rank_by_trend = 8501 // removed
	// cre_rank_by_trend_response = 8502 // removed
	cre_item_vote_summary = 8503
	cre_item_vote_summary_response = 8504
	// cre_rank_by_vote = 8505 // removed
	// cre_rank_by_vote_response = 8506 // removed
	cre_update_user_published_item_vote = 8507
	cre_update_user_published_item_vote_response = 8508
	cre_get_user_published_item_vote_details = 8509
	cre_get_user_published_item_vote_details_response = 8510
	cre_enumerate_published_files = 8511
	cre_enumerate_published_files_response = 8512
	cre_published_file_vote_added = 8513

	// secrets_base = 8600
	secrets_request_credential_pair = 8600
	secrets_credential_pair_response = 8601
	// secrets_request_server_identity = 8602 // removed
	// secrets_server_identity_response = 8603 // removed
	// secrets_update_server_identities = 8604 // removed

	// box_monitor_base = 8700
	box_monitor_report_request = 8700
	box_monitor_report_response = 8701

	// logsink_base = 8800
	logsink_write_report = 8800

	// pics_base = 8900
	client_pics_changes_since_request = 8901
	client_pics_changes_since_response = 8902
	client_pics_product_info_request = 8903
	client_pics_product_info_response = 8904
	client_pics_access_token_request = 8905
	client_pics_access_token_response = 8906

	// worker_process = 9000
	worker_process_ping_request = 9000
	worker_process_ping_response = 9001
	worker_process_shutdown = 9002

	// drm_worker_process = 9100
	drm_worker_process_drm_and_sign = 9100
	drm_worker_process_drm_and_sign_response = 9101
	drm_worker_process_steamworks_info_request = 9102
	drm_worker_process_steamworks_info_response = 9103
	drm_worker_process_install_drmdll_request = 9104
	drm_worker_process_install_drmdll_response = 9105
	drm_worker_process_secret_id_string_request = 9106
	drm_worker_process_secret_id_string_response = 9107
	// drm_worker_process_get_drm_guids_from_file_request = 9108 // removed
	// drm_worker_process_get_drm_guids_from_file_response = 9109 // removed
	drm_worker_process_install_processed_files_request = 9110
	drm_worker_process_install_processed_files_response = 9111
	drm_worker_process_examine_blob_request = 9112
	drm_worker_process_examine_blob_response = 9113
	drm_worker_process_describe_secret_request = 9114
	drm_worker_process_describe_secret_response = 9115
	drm_worker_process_backfill_original_request = 9116
	drm_worker_process_backfill_original_response = 9117
	drm_worker_process_validate_drmdll_request = 9118
	drm_worker_process_validate_drmdll_response = 9119
	drm_worker_process_validate_file_request = 9120
	drm_worker_process_validate_file_response = 9121
	drm_worker_process_split_and_install_request = 9122
	drm_worker_process_split_and_install_response = 9123
	drm_worker_process_get_blob_request = 9124
	drm_worker_process_get_blob_response = 9125
	drm_worker_process_evaluate_crash_request = 9126
	drm_worker_process_evaluate_crash_response = 9127
	drm_worker_process_analyze_file_request = 9128
	drm_worker_process_analyze_file_response = 9129
	drm_worker_process_unpack_blob_request = 9130
	drm_worker_process_unpack_blob_response = 9131
	drm_worker_process_install_all_request = 9132
	drm_worker_process_install_all_response = 9133

	// test_worker_process = 9200
	test_worker_process_load_unload_module_request = 9200
	test_worker_process_load_unload_module_response = 9201
	test_worker_process_service_module_call_request = 9202
	test_worker_process_service_module_call_response = 9203

	// quest_server_base = 9300

	client_get_emoticon_list = 9330
	client_emoticon_list = 9331

	// client_shared_library_base = 9400 // removed "renamed to SLCBase"
	// slc_base = 9400
	slc_user_session_status = 9400
	slc_request_user_session_status = 9401
	slc_shared_licenses_lock_status = 9402
	// client_shared_licenses_lock_status = 9403 // removed
	// client_shared_licenses_stop_playing = 9404 // removed
	client_shared_library_lock_status = 9405
	client_shared_library_stop_playing = 9406
	slc_owner_library_changed = 9407
	slc_shared_library_changed = 9408

	remote_client_base = 9500
	// remote_client_auth = 9500 // obsolete
	// remote_client_auth_response = 9501 // obsolete
	remote_client_app_status = 9502
	remote_client_start_stream = 9503
	remote_client_start_stream_response = 9504
	remote_client_ping = 9505
	remote_client_ping_response = 9506
	client_unlock_streaming = 9507
	client_unlock_streaming_response = 9508
	remote_client_accept_eula = 9509
	remote_client_get_controller_config = 9510
	// remote_client_get_controller_config_resposne = 9511 // obsolete "renamed to RemoteClientGetControllerConfigResponse"
	remote_client_get_controller_config_response = 9511
	remote_client_streaming_enabled = 9512
	client_unlock_hevc = 9513
	client_unlock_hevc_response = 9514
	remote_client_status_request = 9515
	remote_client_status_response = 9516

	// client_concurrent_sessions_base = 9600
	client_playing_session_state = 9600
	client_kick_playing_session = 9601

	// client_broadcast_base = 9700
	client_broadcast_init = 9700
	client_broadcast_frames = 9701
	client_broadcast_disconnect = 9702
	client_broadcast_screenshot = 9703
	client_broadcast_upload_config = 9704

	// base_client3 = 9800
	client_voice_call_pre_authorize = 9800
	client_voice_call_pre_authorize_response = 9801
	client_server_timestamp_request = 9802
	client_server_timestamp_response = 9803

	// client_lanp2_p_base = 9900
	client_lanp2_p_request_chunk = 9900
	client_lanp2_p_request_chunk_response = 9901
	client_lanp2_p_max = 9999

	// base_watchdog_server = 10000
	notify_watchdog = 10000

	// client_site_license_base = 10100
	client_site_license_site_info_notification = 10100
	client_site_license_checkout = 10101
	client_site_license_checkout_response = 10102
	client_site_license_get_available_seats = 10103
	client_site_license_get_available_seats_response = 10104
	client_site_license_get_content_cache_info = 10105
	client_site_license_get_content_cache_info_response = 10106

	// base_chat_server = 12000
	chat_server_get_pending_notification_count = 12000
	chat_server_get_pending_notification_count_response = 12001

	// base_secret_server = 12100
	server_secret_changed = 12100
}

pub fn (m Msg) make_proto() u32 {
	return msg_make_proto(m)
}

const (
	proto_mask = 0x80000000
)

fn msg_is_proto(msg u32) bool {
	return msg & proto_mask == proto_mask
}

fn msg_make_proto(msg Msg) u32 {
	return u32(msg) | proto_mask
}

fn raw_msg(msg u32) Msg {
	return Msg(msg & ~proto_mask)
}