module vapor

struct SteamFriends {
}

pub fn (mut s SteamFriends) initialise() ? {
	
}

pub fn (mut s SteamFriends) handle_msg(mut m Message) ? {

}